module constant0 (
    output y
    );
    assign y = 1'b0;
    
endmodule
